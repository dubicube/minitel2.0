--|==========================================================================|--
--|  ____        _    _  _              _                                    |--
--| |    \  _ _ | |_ |_|| |_  ___  ___ | |_                                  |--
--| |  |  || | || . || ||  _|| -_||  _||   |                                 |--
--| |____/ |___||___||_||_|  |___||___||_|_|                                 |--
--|                                                                          |--
--|==========================================================================|--
--| Module name: ascii_converter                                             |--
--| Description: Converts keyboard matrix data to ascii characters           |--
--|                                                                          |--
--|==========================================================================|--
--| 31/12/2020 | Creation                                                    |--
--|            |                                                             |--
--|==========================================================================|--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;
--library UNISIM;
--use UNISIM.VComponents.all;

entity ascii_converter is
Port (
   CLK : in std_logic;

   -- Keyboard input
   KEY_UPDATE : in std_logic;
   KEY_REG    : in std_logic_vector(63 downto 0);

   -- ASCII output
   CHAR_VALID : out std_logic;
   CHAR_DATA  : out std_logic_vector(7 downto 0)
);
end ascii_converter;

architecture Behavioral of ascii_converter is
   --|=======================================================================|--
   --| Internal signals
   --|=======================================================================|--

   -- Just an ASCII table, but special (generated from table.py script)
   type t_MEMORY_16 is array (0 to 1023) of integer range 0 to 511;
   -- Integers because we cant express 9 bits values in hexadecimal in VHDL (I didnt found the way to do it on stack overflow...)
   constant c_ASCII_TABLE : t_MEMORY_16 := (
      283, 347, 305, 321, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 283, 347, 305, 322, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 283, 347, 305, 324, 0, 0, 0, 0, 283, 347, 305, 323, 0, 0, 0, 0, 269, 0, 0, 0, 0, 0, 0, 0,
      372, 0, 0, 0, 0, 0, 0, 0, 357, 0, 0, 0, 0, 0, 0, 0, 370, 0, 0, 0, 0, 0, 0, 0, 377, 0, 0, 0, 0, 0, 0, 0,
      315, 0, 0, 0, 0, 0, 0, 0, 301, 0, 0, 0, 0, 0, 0, 0, 314, 0, 0, 0, 0, 0, 0, 0, 319, 0, 0, 0, 0, 0, 0, 0,
      359, 0, 0, 0, 0, 0, 0, 0, 356, 0, 0, 0, 0, 0, 0, 0, 358, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 0, 0, 0, 0, 0,
      298, 0, 0, 0, 0, 0, 0, 0, 311, 0, 0, 0, 0, 0, 0, 0, 308, 0, 0, 0, 0, 0, 0, 0, 305, 0, 0, 0, 0, 0, 0, 0,
      302, 0, 0, 0, 0, 0, 0, 0, 283, 0, 0, 0, 0, 0, 0, 0, 300, 0, 0, 0, 0, 0, 0, 0, 295, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      354, 0, 0, 0, 0, 0, 0, 0, 355, 0, 0, 0, 0, 0, 0, 0, 374, 0, 0, 0, 0, 0, 0, 0, 366, 0, 0, 0, 0, 0, 0, 0,
      304, 0, 0, 0, 0, 0, 0, 0, 312, 0, 0, 0, 0, 0, 0, 0, 309, 0, 0, 0, 0, 0, 0, 0, 306, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 378, 0, 0, 0, 0, 0, 0, 0, 353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      373, 0, 0, 0, 0, 0, 0, 0, 361, 0, 0, 0, 0, 0, 0, 0, 367, 0, 0, 0, 0, 0, 0, 0, 368, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 371, 0, 0, 0, 0, 0, 0, 0, 369, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      362, 0, 0, 0, 0, 0, 0, 0, 363, 0, 0, 0, 0, 0, 0, 0, 364, 0, 0, 0, 0, 0, 0, 0, 365, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 376, 0, 0, 0, 0, 0, 0, 0, 375, 0, 0, 0, 0, 0, 0, 0, 288, 0, 0, 0, 0, 0, 0, 0,
      291, 0, 0, 0, 0, 0, 0, 0, 313, 0, 0, 0, 0, 0, 0, 0, 310, 0, 0, 0, 0, 0, 0, 0, 307, 0, 0, 0, 0, 0, 0, 0,
      283, 347, 305, 321, 0, 0, 0, 0, 501, 0, 0, 0, 0, 0, 0, 0, 348, 0, 0, 0, 0, 0, 0, 0, 283, 347, 305, 322, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 283, 347, 305, 324, 0, 0, 0, 0, 283, 347, 305, 323, 0, 0, 0, 0, 266, 0, 0, 0, 0, 0, 0, 0,
      340, 0, 0, 0, 0, 0, 0, 0, 325, 0, 0, 0, 0, 0, 0, 0, 338, 0, 0, 0, 0, 0, 0, 0, 345, 0, 0, 0, 0, 0, 0, 0,
      299, 0, 0, 0, 0, 0, 0, 0, 317, 0, 0, 0, 0, 0, 0, 0, 298, 0, 0, 0, 0, 0, 0, 0, 303, 0, 0, 0, 0, 0, 0, 0,
      327, 0, 0, 0, 0, 0, 0, 0, 324, 0, 0, 0, 0, 0, 0, 0, 326, 0, 0, 0, 0, 0, 0, 0, 328, 0, 0, 0, 0, 0, 0, 0,
      347, 0, 0, 0, 0, 0, 0, 0, 295, 0, 0, 0, 0, 0, 0, 0, 292, 0, 0, 0, 0, 0, 0, 0, 289, 0, 0, 0, 0, 0, 0, 0,
      318, 0, 0, 0, 0, 0, 0, 0, 283, 0, 0, 0, 0, 0, 0, 0, 316, 0, 0, 0, 0, 0, 0, 0, 320, 0, 0, 0, 0, 0, 0, 0,
      352, 0, 0, 0, 0, 0, 0, 0, 495, 0, 0, 0, 0, 0, 0, 0, 381, 0, 0, 0, 0, 0, 0, 0, 379, 0, 0, 0, 0, 0, 0, 0,
      322, 0, 0, 0, 0, 0, 0, 0, 323, 0, 0, 0, 0, 0, 0, 0, 342, 0, 0, 0, 0, 0, 0, 0, 334, 0, 0, 0, 0, 0, 0, 0,
      424, 0, 0, 0, 0, 0, 0, 0, 296, 0, 0, 0, 0, 0, 0, 0, 293, 0, 0, 0, 0, 0, 0, 0, 290, 0, 0, 0, 0, 0, 0, 0,
      505, 0, 0, 0, 0, 0, 0, 0, 346, 0, 0, 0, 0, 0, 0, 0, 321, 0, 0, 0, 0, 0, 0, 0, 350, 0, 0, 0, 0, 0, 0, 0,
      341, 0, 0, 0, 0, 0, 0, 0, 329, 0, 0, 0, 0, 0, 0, 0, 335, 0, 0, 0, 0, 0, 0, 0, 336, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 339, 0, 0, 0, 0, 0, 0, 0, 337, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      330, 0, 0, 0, 0, 0, 0, 0, 331, 0, 0, 0, 0, 0, 0, 0, 332, 0, 0, 0, 0, 0, 0, 0, 333, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 344, 0, 0, 0, 0, 0, 0, 0, 343, 0, 0, 0, 0, 0, 0, 0, 288, 0, 0, 0, 0, 0, 0, 0,
      349, 0, 0, 0, 0, 0, 0, 0, 297, 0, 0, 0, 0, 0, 0, 0, 294, 0, 0, 0, 0, 0, 0, 0, 291, 0, 0, 0, 0, 0, 0, 0
   );

   signal s_KEY_REG_d1 : std_logic_vector(63 downto 0) := (others => '1');
   -- signal s_KEY_REG_d2 : std_logic_vector(63 downto 0) := (others => '1');
   signal s_KEY_UPDATE : std_logic := '0';

   signal s_step        : unsigned(5 downto 0) := (others => '0');
   signal s_step_i      : integer range 0 to 63;
   signal s_char_num    : unsigned(2 downto 0) := (others => '0');
   signal s_table_index : unsigned(1 downto 0);

   signal s_sweep_finished : std_logic;

   signal s_rom_addr   : unsigned(9 downto 0);
   signal s_rom_addr_i : integer range 0 to (2**10)-1;
   signal s_rom_data   : std_logic_vector(8 downto 0);

   signal s_CHAR_VALID : std_logic := '0';

begin

   s_table_index(0) <= not KEY_REG(4);
   s_table_index(1) <= '0';

   --|=======================================================================|--
   --| Char output
   --|=======================================================================|--
   CHAR_DATA  <= s_rom_data(7 downto 0);
   CHAR_VALID <= s_CHAR_VALID and s_rom_data(8);
   process(CLK) begin
      if rising_edge(CLK) then
         if (s_sweep_finished = '0' and KEY_REG(s_step_i) = '0' and s_KEY_REG_d1(s_step_i) = '1') then
            s_CHAR_VALID <= '1';
         else
            s_CHAR_VALID <= '0';
         end if;
      end if;
   end process;
   s_step_i <= to_integer(s_step);

   --|=======================================================================|--
   --| Counters
   --|=======================================================================|--
   process(CLK) begin
      if rising_edge(CLK) then
         if (s_char_num /= "111" or s_step /= "111111" or s_KEY_UPDATE = '1') then
            s_char_num <= s_char_num + 1;
            if (s_char_num = "111") then
               s_step <= s_step + 1;
            end if;
            s_sweep_finished <= '0';
         else
            s_sweep_finished <= '1';
         end if;
      end if;
   end process;

   --|=======================================================================|--
   --| ROM
   --|=======================================================================|--
   s_rom_addr_i <= to_integer(s_rom_addr);
   s_rom_addr <= s_table_index(0 downto 0) & s_step & s_char_num;
   process(CLK) begin
      if rising_edge(CLK) then
         s_rom_data <= std_logic_vector(to_unsigned(c_ASCII_TABLE(s_rom_addr_i), 9));
      end if;
   end process;

   --|=======================================================================|--
   --| Keyboard input
   --|=======================================================================|--
   process(CLK) begin
      if rising_edge(CLK) then
         if (s_sweep_finished = '0' and s_char_num = "111" and s_step = "111111") then
            s_KEY_REG_d1 <= KEY_REG;
            -- s_KEY_REG_d2 <= s_KEY_REG_d1;
         end if;
         s_KEY_UPDATE <= KEY_UPDATE;
      end if;
   end process;

end Behavioral;
