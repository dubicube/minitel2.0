--|==========================================================================|--
--|  ____        _    _  _              _                                    |--
--| |    \  _ _ | |_ |_|| |_  ___  ___ | |_                                  |--
--| |  |  || | || . || ||  _|| -_||  _||   |                                 |--
--| |____/ |___||___||_||_|  |___||___||_|_|                                 |--
--|                                                                          |--
--|==========================================================================|--
--| Module name: ascii_converter                                             |--
--| Description: Converts keyboard matrix data to ascii characters           |--
--|                                                                          |--
--|==========================================================================|--
--| 31/12/2020 | Creation                                                    |--
--|            |                                                             |--
--|==========================================================================|--

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;
--library UNISIM;
--use UNISIM.VComponents.all;

entity ascii_converter is
Port (
   CLK : in std_logic;

   -- Keyboard input
   KEY_UPDATE : in std_logic;
   KEY_REG    : in std_logic_vector(63 downto 0)

   -- ASCII output
   CHAR_READY : in  std_logic;
   CHAR_VALID : out std_logic;
   CHAR_DATA  : out std_logic_vector(7 downto 0)
);
end ascii_converter;

architecture Behavioral of ascii_converter is
   --|=======================================================================|--
   --| Internal signals
   --|=======================================================================|--

   -- Just an ASCII table, but special (generated from table.py script)
   type t_MEMORY_16 is array (0 to 1023) of integer range 0 to 511;
   -- Integers because we cant express 9 bits values in hexadecimal in VHDL (I didnt found the way to do it on stack overflow...)
   constant c_ASCII_TABLE : t_MEMORY_16 := (
      27, 91, 49, 321, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 27, 91, 49, 322, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 27, 91, 49, 324, 256, 256, 256, 256, 27, 91, 49, 323, 256, 256, 256, 256, 269, 256, 256, 256, 256, 256, 256, 256,
      372, 256, 256, 256, 256, 256, 256, 256, 357, 256, 256, 256, 256, 256, 256, 256, 370, 256, 256, 256, 256, 256, 256, 256, 377, 256, 256, 256, 256, 256, 256, 256,
      315, 256, 256, 256, 256, 256, 256, 256, 301, 256, 256, 256, 256, 256, 256, 256, 314, 256, 256, 256, 256, 256, 256, 256, 319, 256, 256, 256, 256, 256, 256, 256,
      359, 256, 256, 256, 256, 256, 256, 256, 356, 256, 256, 256, 256, 256, 256, 256, 358, 256, 256, 256, 256, 256, 256, 256, 360, 256, 256, 256, 256, 256, 256, 256,
      298, 256, 256, 256, 256, 256, 256, 256, 311, 256, 256, 256, 256, 256, 256, 256, 308, 256, 256, 256, 256, 256, 256, 256, 305, 256, 256, 256, 256, 256, 256, 256,
      302, 256, 256, 256, 256, 256, 256, 256, 283, 256, 256, 256, 256, 256, 256, 256, 300, 256, 256, 256, 256, 256, 256, 256, 295, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256,
      354, 256, 256, 256, 256, 256, 256, 256, 355, 256, 256, 256, 256, 256, 256, 256, 374, 256, 256, 256, 256, 256, 256, 256, 366, 256, 256, 256, 256, 256, 256, 256,
      304, 256, 256, 256, 256, 256, 256, 256, 312, 256, 256, 256, 256, 256, 256, 256, 341, 256, 256, 256, 256, 256, 256, 256, 306, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 378, 256, 256, 256, 256, 256, 256, 256, 353, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256,
      373, 256, 256, 256, 256, 256, 256, 256, 361, 256, 256, 256, 256, 256, 256, 256, 367, 256, 256, 256, 256, 256, 256, 256, 368, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 371, 256, 256, 256, 256, 256, 256, 256, 369, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256,
      362, 256, 256, 256, 256, 256, 256, 256, 363, 256, 256, 256, 256, 256, 256, 256, 364, 256, 256, 256, 256, 256, 256, 256, 365, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 376, 256, 256, 256, 256, 256, 256, 256, 375, 256, 256, 256, 256, 256, 256, 256, 288, 256, 256, 256, 256, 256, 256, 256,
      291, 256, 256, 256, 256, 256, 256, 256, 313, 256, 256, 256, 256, 256, 256, 256, 310, 256, 256, 256, 256, 256, 256, 256, 307, 256, 256, 256, 256, 256, 256, 256,
      27, 91, 49, 321, 256, 256, 256, 256, 501, 256, 256, 256, 256, 256, 256, 256, 348, 256, 256, 256, 256, 256, 256, 256, 27, 91, 49, 322, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 27, 91, 49, 324, 256, 256, 256, 256, 27, 91, 49, 323, 256, 256, 256, 256, 266, 256, 256, 256, 256, 256, 256, 256,
      340, 256, 256, 256, 256, 256, 256, 256, 325, 256, 256, 256, 256, 256, 256, 256, 338, 256, 256, 256, 256, 256, 256, 256, 345, 256, 256, 256, 256, 256, 256, 256,
      299, 256, 256, 256, 256, 256, 256, 256, 317, 256, 256, 256, 256, 256, 256, 256, 298, 256, 256, 256, 256, 256, 256, 256, 303, 256, 256, 256, 256, 256, 256, 256,
      327, 256, 256, 256, 256, 256, 256, 256, 324, 256, 256, 256, 256, 256, 256, 256, 326, 256, 256, 256, 256, 256, 256, 256, 328, 256, 256, 256, 256, 256, 256, 256,
      347, 256, 256, 256, 256, 256, 256, 256, 295, 256, 256, 256, 256, 256, 256, 256, 292, 256, 256, 256, 256, 256, 256, 256, 289, 256, 256, 256, 256, 256, 256, 256,
      318, 256, 256, 256, 256, 256, 256, 256, 283, 256, 256, 256, 256, 256, 256, 256, 316, 256, 256, 256, 256, 256, 256, 256, 320, 256, 256, 256, 256, 256, 256, 256,
      352, 256, 256, 256, 256, 256, 256, 256, 495, 256, 256, 256, 256, 256, 256, 256, 381, 256, 256, 256, 256, 256, 256, 256, 379, 256, 256, 256, 256, 256, 256, 256,
      322, 256, 256, 256, 256, 256, 256, 256, 323, 256, 256, 256, 256, 256, 256, 256, 342, 256, 256, 256, 256, 256, 256, 256, 334, 256, 256, 256, 256, 256, 256, 256,
      424, 256, 256, 256, 256, 256, 256, 256, 296, 256, 256, 256, 256, 256, 256, 256, 293, 256, 256, 256, 256, 256, 256, 256, 290, 256, 256, 256, 256, 256, 256, 256,
      505, 256, 256, 256, 256, 256, 256, 256, 346, 256, 256, 256, 256, 256, 256, 256, 321, 256, 256, 256, 256, 256, 256, 256, 350, 256, 256, 256, 256, 256, 256, 256,
      341, 256, 256, 256, 256, 256, 256, 256, 329, 256, 256, 256, 256, 256, 256, 256, 335, 256, 256, 256, 256, 256, 256, 256, 336, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 339, 256, 256, 256, 256, 256, 256, 256, 337, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256, 256,
      330, 256, 256, 256, 256, 256, 256, 256, 331, 256, 256, 256, 256, 256, 256, 256, 332, 256, 256, 256, 256, 256, 256, 256, 333, 256, 256, 256, 256, 256, 256, 256,
      256, 256, 256, 256, 256, 256, 256, 256, 344, 256, 256, 256, 256, 256, 256, 256, 343, 256, 256, 256, 256, 256, 256, 256, 288, 256, 256, 256, 256, 256, 256, 256,
      349, 256, 256, 256, 256, 256, 256, 256, 297, 256, 256, 256, 256, 256, 256, 256, 294, 256, 256, 256, 256, 256, 256, 256, 291, 256, 256, 256, 256, 256, 256, 256
   );

   signal s_KEY_REG    : std_logic_vector(63 downto 0) := (others => '1');
   signal s_KEY_UPDATE : std_logic := '0';

   signal s_step        : unsigned(5 downto 0) := (others => '0');
   signal s_char_num    : unsigned(2 downto 0) := (others => '0');
   signal s_table_index : unsigned(1 downto 0) := (others => '0');

   signal s_next_step : std_logic;
   signal s_next_char : std_logic;

   signal s_rom_addr : std_logic_vector(9 downto 0);
   signal s_rom_data : std_logic_vector(8 downto 0);

begin

   s_rom_addr <= s_table_index(0 downto 0) & s_step & s_char_num;

   s_next_step <= '1' when KEY_UPDATE = '1' else '0';
   s_next_char <= '1' when s_rom_data(8)='0' else '0';


   --|=======================================================================|--
   --|
   --|=======================================================================|--
   process(CLK) begin
      if rising_edge(CLK) then
         if (s_next_step = '1') then
            s_step <= s_step + 1;
            s_char_num <= (others => '0');
         end if;
      end if;
   end process;

   --|=======================================================================|--
   --| ROM
   --|=======================================================================|--
   process(CLK) begin
      if rising_edge(CLK) then
         s_rom_data <= c_ASCII_TABLE(s_rom_addr);
      end if;
   end process;

   --|=======================================================================|--
   --| Keyboard input
   --|=======================================================================|--
   process(CLK) begin
      if rising_edge(CLK) then
         if (KEY_UPDATE = '1') then
            s_KEY_REG <= KEY_REG;
         end if;
         s_KEY_UPDATE <= KEY_UPDATE;
      end if;
   end process;

end Behavioral;
